module Seven_segment_Decoder(input [3:0] a ,
output [6:0] c);

assign c= (a=== 4'b0000)?  7'b1000_000  :
 (a=== 4'b0001)? 7'b1111_001:
 (a=== 4'b0010)? 7'b0100_100:
 (a=== 4'b0011)? 7'b0110_000:
 (a=== 4'b0100)? 7'b0011_001:
 (a=== 4'b0101)? 7'b0010_010:
 (a=== 4'b0110)? 7'b0000_010:
 (a=== 4'b0111)? 7'b1111_000:
 (a=== 4'b1000)? 7'b0000_000:
 (a=== 4'b1001)? 7'b0010_000:
7'b1000_000;

endmodule